-- nios_hps_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_hps_system is
	port (
		clk_clk                            : in    std_logic                     := '0';             --                     clk.clk
		hps_0_ddr_mem_a                    : out   std_logic_vector(14 downto 0);                    --               hps_0_ddr.mem_a
		hps_0_ddr_mem_ba                   : out   std_logic_vector(2 downto 0);                     --                        .mem_ba
		hps_0_ddr_mem_ck                   : out   std_logic;                                        --                        .mem_ck
		hps_0_ddr_mem_ck_n                 : out   std_logic;                                        --                        .mem_ck_n
		hps_0_ddr_mem_cke                  : out   std_logic;                                        --                        .mem_cke
		hps_0_ddr_mem_cs_n                 : out   std_logic;                                        --                        .mem_cs_n
		hps_0_ddr_mem_ras_n                : out   std_logic;                                        --                        .mem_ras_n
		hps_0_ddr_mem_cas_n                : out   std_logic;                                        --                        .mem_cas_n
		hps_0_ddr_mem_we_n                 : out   std_logic;                                        --                        .mem_we_n
		hps_0_ddr_mem_reset_n              : out   std_logic;                                        --                        .mem_reset_n
		hps_0_ddr_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => '0'); --                        .mem_dq
		hps_0_ddr_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs
		hps_0_ddr_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs_n
		hps_0_ddr_mem_odt                  : out   std_logic;                                        --                        .mem_odt
		hps_0_ddr_mem_dm                   : out   std_logic_vector(3 downto 0);                     --                        .mem_dm
		hps_0_ddr_oct_rzqin                : in    std_logic                     := '0';             --                        .oct_rzqin
		hps_0_h2f_loan_io_in               : out   std_logic_vector(66 downto 0);                    --       hps_0_h2f_loan_io.in
		hps_0_h2f_loan_io_out              : in    std_logic_vector(66 downto 0) := (others => '0'); --                        .out
		hps_0_h2f_loan_io_oe               : in    std_logic_vector(66 downto 0) := (others => '0'); --                        .oe
		hps_0_io_hps_io_sdio_inst_CMD      : inout std_logic                     := '0';             --                hps_0_io.hps_io_sdio_inst_CMD
		hps_0_io_hps_io_sdio_inst_D0       : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D0
		hps_0_io_hps_io_sdio_inst_D1       : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D1
		hps_0_io_hps_io_sdio_inst_CLK      : out   std_logic;                                        --                        .hps_io_sdio_inst_CLK
		hps_0_io_hps_io_sdio_inst_D2       : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D2
		hps_0_io_hps_io_sdio_inst_D3       : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D3
		hps_0_io_hps_io_gpio_inst_LOANIO49 : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_LOANIO49
		hps_0_io_hps_io_gpio_inst_LOANIO50 : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_LOANIO50
		hps_0_io_hps_io_gpio_inst_LOANIO55 : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_LOANIO55
		hps_0_io_hps_io_gpio_inst_LOANIO56 : inout std_logic                     := '0';             --                        .hps_io_gpio_inst_LOANIO56
		i2c_peripheral_sda_in              : in    std_logic                     := '0';             --          i2c_peripheral.sda_in
		i2c_peripheral_scl_in              : in    std_logic                     := '0';             --                        .scl_in
		i2c_peripheral_sda_oe              : out   std_logic;                                        --                        .sda_oe
		i2c_peripheral_scl_oe              : out   std_logic;                                        --                        .scl_oe
		nios_7seg_export                   : out   std_logic_vector(23 downto 0);                    --               nios_7seg.export
		nios_buttons_export                : in    std_logic_vector(3 downto 0)  := (others => '0'); --            nios_buttons.export
		nios_header_conn_in_port           : in    std_logic_vector(31 downto 0) := (others => '0'); --        nios_header_conn.in_port
		nios_header_conn_out_port          : out   std_logic_vector(31 downto 0);                    --                        .out_port
		nios_i2cclk_export                 : out   std_logic;                                        --             nios_i2cclk.export
		nios_i2cdat_in_port                : in    std_logic                     := '0';             --             nios_i2cdat.in_port
		nios_i2cdat_out_port               : out   std_logic;                                        --                        .out_port
		nios_i2crw_export                  : out   std_logic;                                        --              nios_i2crw.export
		nios_leds_export                   : out   std_logic_vector(9 downto 0);                     --               nios_leds.export
		nios_oscdivisor_export             : out   std_logic_vector(15 downto 0);                    --         nios_oscdivisor.export
		nios_switches_export               : in    std_logic_vector(9 downto 0)  := (others => '0'); --           nios_switches.export
		nios_uartrx_export                 : in    std_logic                     := '0';             --             nios_uartrx.export
		nios_uarttx_export                 : out   std_logic;                                        --             nios_uarttx.export
		pll_0_sdram_clk                    : out   std_logic;                                        --             pll_0_sdram.clk
		pll_1_108_clk                      : out   std_logic;                                        --               pll_1_108.clk
		pll_1_144_clk                      : out   std_logic;                                        --               pll_1_144.clk
		pll_1_162_clk                      : out   std_logic;                                        --               pll_1_162.clk
		pll_1_65_clk                       : out   std_logic;                                        --                pll_1_65.clk
		pll_1_86_clk                       : out   std_logic;                                        --                pll_1_86.clk
		reset_reset_n                      : in    std_logic                     := '0';             --                   reset.reset_n
		sdram_controller_0_wire_addr       : out   std_logic_vector(12 downto 0);                    -- sdram_controller_0_wire.addr
		sdram_controller_0_wire_ba         : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_controller_0_wire_cas_n      : out   std_logic;                                        --                        .cas_n
		sdram_controller_0_wire_cke        : out   std_logic;                                        --                        .cke
		sdram_controller_0_wire_cs_n       : out   std_logic;                                        --                        .cs_n
		sdram_controller_0_wire_dq         : inout std_logic_vector(15 downto 0) := (others => '0'); --                        .dq
		sdram_controller_0_wire_dqm        : out   std_logic_vector(1 downto 0);                     --                        .dqm
		sdram_controller_0_wire_ras_n      : out   std_logic;                                        --                        .ras_n
		sdram_controller_0_wire_we_n       : out   std_logic;                                        --                        .we_n
		spi_peripheral_MISO                : in    std_logic                     := '0';             --          spi_peripheral.MISO
		spi_peripheral_MOSI                : out   std_logic;                                        --                        .MOSI
		spi_peripheral_SCLK                : out   std_logic;                                        --                        .SCLK
		spi_peripheral_SS_n                : out   std_logic;                                        --                        .SS_n
		uart_peripheral_rxd                : in    std_logic                     := '0';             --         uart_peripheral.rxd
		uart_peripheral_txd                : out   std_logic                                         --                        .txd
	);
end entity nios_hps_system;

architecture rtl of nios_hps_system is
	component nios_hps_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_loan_in               : out   std_logic_vector(66 downto 0);                    -- in
			h2f_loan_out              : in    std_logic_vector(66 downto 0) := (others => 'X'); -- out
			h2f_loan_oe               : in    std_logic_vector(66 downto 0) := (others => 'X'); -- oe
			mem_a                     : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                    : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                    : out   std_logic;                                        -- mem_ck
			mem_ck_n                  : out   std_logic;                                        -- mem_ck_n
			mem_cke                   : out   std_logic;                                        -- mem_cke
			mem_cs_n                  : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                 : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                 : out   std_logic;                                        -- mem_cas_n
			mem_we_n                  : out   std_logic;                                        -- mem_we_n
			mem_reset_n               : out   std_logic;                                        -- mem_reset_n
			mem_dq                    : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                   : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                 : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                   : out   std_logic;                                        -- mem_odt
			mem_dm                    : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                 : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_sdio_inst_CMD      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0       : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1       : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK      : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2       : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3       : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_gpio_inst_LOANIO49 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO49
			hps_io_gpio_inst_LOANIO50 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO50
			hps_io_gpio_inst_LOANIO55 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO55
			hps_io_gpio_inst_LOANIO56 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO56
			h2f_rst_n                 : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk            : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID               : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR             : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN              : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE             : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST            : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK             : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE            : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT             : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID            : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY            : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID                : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA              : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB              : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST              : out   std_logic;                                        -- wlast
			h2f_lw_WVALID             : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY             : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID                : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID             : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY             : out   std_logic;                                        -- bready
			h2f_lw_ARID               : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR             : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN              : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE             : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST            : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK             : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE            : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT             : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID            : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY            : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID                : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA              : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST              : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID             : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY             : out   std_logic                                         -- rready
		);
	end component nios_hps_system_hps_0;

	component altera_avalon_i2c is
		generic (
			USE_AV_ST       : integer := 0;
			FIFO_DEPTH      : integer := 4;
			FIFO_DEPTH_LOG2 : integer := 2
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			rst_n     : in  std_logic                     := 'X';             -- reset_n
			intr      : out std_logic;                                        -- irq
			addr      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			sda_in    : in  std_logic                     := 'X';             -- sda_in
			scl_in    : in  std_logic                     := 'X';             -- scl_in
			sda_oe    : out std_logic;                                        -- sda_oe
			scl_oe    : out std_logic;                                        -- scl_oe
			src_data  : out std_logic_vector(7 downto 0);                     -- data
			src_valid : out std_logic;                                        -- valid
			src_ready : in  std_logic                     := 'X';             -- ready
			snk_data  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			snk_valid : in  std_logic                     := 'X';             -- valid
			snk_ready : out std_logic                                         -- ready
		);
	end component altera_avalon_i2c;

	component nios_hps_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_hps_system_jtag_uart_0;

	component nios_hps_system_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(27 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios_hps_system_nios2_qsys_0;

	component nios_hps_system_nios_7seg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(23 downto 0)                     -- export
		);
	end component nios_hps_system_nios_7seg;

	component nios_hps_system_nios_buttons is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component nios_hps_system_nios_buttons;

	component nios_hps_system_nios_header_conn is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component nios_hps_system_nios_header_conn;

	component nios_hps_system_nios_i2cclk is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_hps_system_nios_i2cclk;

	component nios_hps_system_nios_i2cdat is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			out_port   : out std_logic                                         -- export
		);
	end component nios_hps_system_nios_i2cdat;

	component nios_hps_system_nios_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component nios_hps_system_nios_leds;

	component nios_hps_system_nios_oscdivisor is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component nios_hps_system_nios_oscdivisor;

	component nios_hps_system_nios_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component nios_hps_system_nios_switches;

	component nios_hps_system_nios_uartrx is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component nios_hps_system_nios_uartrx;

	component nios_hps_system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component nios_hps_system_pll_0;

	component nios_hps_system_pll_1 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			outclk_3 : out std_logic;        -- clk
			outclk_4 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component nios_hps_system_pll_1;

	component nios_hps_system_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_hps_system_sdram_controller_0;

	component nios_hps_system_spi_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_hps_system_spi_0;

	component nios_hps_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_hps_system_sysid_qsys_0;

	component nios_hps_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_hps_system_timer_0;

	component nios_hps_system_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component nios_hps_system_uart_0;

	component nios_hps_system_mm_interconnect_0 is
		port (
			pll_0_outclk0_clk                                : in  std_logic                     := 'X';             -- clk
			pll_0_outclk1_clk                                : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_data_master_address                 : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address          : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			i2c_0_csr_address                                : out std_logic_vector(3 downto 0);                     -- address
			i2c_0_csr_write                                  : out std_logic;                                        -- write
			i2c_0_csr_read                                   : out std_logic;                                        -- read
			i2c_0_csr_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_0_csr_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_address            : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write              : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read               : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect         : out std_logic;                                        -- chipselect
			nios2_qsys_0_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_qsys_0_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_qsys_0_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			nios_7seg_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			nios_7seg_s1_write                               : out std_logic;                                        -- write
			nios_7seg_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_7seg_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			nios_7seg_s1_chipselect                          : out std_logic;                                        -- chipselect
			nios_buttons_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			nios_buttons_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_header_conn_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			nios_header_conn_s1_write                        : out std_logic;                                        -- write
			nios_header_conn_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_header_conn_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			nios_header_conn_s1_chipselect                   : out std_logic;                                        -- chipselect
			nios_i2cclk_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			nios_i2cclk_s1_write                             : out std_logic;                                        -- write
			nios_i2cclk_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_i2cclk_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			nios_i2cclk_s1_chipselect                        : out std_logic;                                        -- chipselect
			nios_i2cdat_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			nios_i2cdat_s1_write                             : out std_logic;                                        -- write
			nios_i2cdat_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_i2cdat_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			nios_i2cdat_s1_chipselect                        : out std_logic;                                        -- chipselect
			nios_i2crw_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			nios_i2crw_s1_write                              : out std_logic;                                        -- write
			nios_i2crw_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_i2crw_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			nios_i2crw_s1_chipselect                         : out std_logic;                                        -- chipselect
			nios_leds_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			nios_leds_s1_write                               : out std_logic;                                        -- write
			nios_leds_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_leds_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			nios_leds_s1_chipselect                          : out std_logic;                                        -- chipselect
			nios_oscdivisor_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nios_oscdivisor_s1_write                         : out std_logic;                                        -- write
			nios_oscdivisor_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_oscdivisor_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nios_oscdivisor_s1_chipselect                    : out std_logic;                                        -- chipselect
			nios_switches_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			nios_switches_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_uartrx_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			nios_uartrx_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_uarttx_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			nios_uarttx_s1_write                             : out std_logic;                                        -- write
			nios_uarttx_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_uarttx_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			nios_uarttx_s1_chipselect                        : out std_logic;                                        -- chipselect
			sdram_controller_0_s1_address                    : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_0_s1_write                      : out std_logic;                                        -- write
			sdram_controller_0_s1_read                       : out std_logic;                                        -- read
			sdram_controller_0_s1_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_0_s1_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_0_s1_byteenable                 : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_0_s1_readdatavalid              : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_0_s1_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			spi_0_spi_control_port_address                   : out std_logic_vector(2 downto 0);                     -- address
			spi_0_spi_control_port_write                     : out std_logic;                                        -- write
			spi_0_spi_control_port_read                      : out std_logic;                                        -- read
			spi_0_spi_control_port_readdata                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_0_spi_control_port_writedata                 : out std_logic_vector(15 downto 0);                    -- writedata
			spi_0_spi_control_port_chipselect                : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                               : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                 : out std_logic;                                        -- write
			timer_0_s1_readdata                              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                             : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                            : out std_logic;                                        -- chipselect
			uart_0_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                                  : out std_logic;                                        -- write
			uart_0_s1_read                                   : out std_logic;                                        -- read
			uart_0_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer                          : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                             : out std_logic                                         -- chipselect
		);
	end component nios_hps_system_mm_interconnect_0;

	component nios_hps_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_hps_system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component nios_hps_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_hps_system_rst_controller;

	component nios_hps_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_hps_system_rst_controller_001;

	signal pll_0_outclk0_clk                                               : std_logic;                     -- pll_0:outclk_0 -> [hps_0:h2f_lw_axi_clk, i2c_0:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, irq_synchronizer_004:receiver_clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, nios_7seg:clk, nios_buttons:clk, nios_header_conn:clk, nios_i2cclk:clk, nios_i2cdat:clk, nios_i2crw:clk, nios_leds:clk, nios_oscdivisor:clk, nios_switches:clk, nios_uartrx:clk, nios_uarttx:clk, rst_controller:clk, spi_0:clk, sysid_qsys_0:clock, timer_0:clk, uart_0:clk]
	signal pll_0_outclk1_clk                                               : std_logic;                     -- pll_0:outclk_1 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, mm_interconnect_0:pll_0_outclk1_clk, nios2_qsys_0:clk, rst_controller_001:clk, sdram_controller_0:clk]
	signal nios2_qsys_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_debugaccess                            : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_address                                : std_logic_vector(27 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal nios2_qsys_0_data_master_read                                   : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_write                                  : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal nios2_qsys_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                         : std_logic_vector(27 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                            : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_i2c_0_csr_readdata                            : std_logic_vector(31 downto 0); -- i2c_0:readdata -> mm_interconnect_0:i2c_0_csr_readdata
	signal mm_interconnect_0_i2c_0_csr_address                             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:i2c_0_csr_address -> i2c_0:addr
	signal mm_interconnect_0_i2c_0_csr_read                                : std_logic;                     -- mm_interconnect_0:i2c_0_csr_read -> i2c_0:read
	signal mm_interconnect_0_i2c_0_csr_write                               : std_logic;                     -- mm_interconnect_0:i2c_0_csr_write -> i2c_0:write
	signal mm_interconnect_0_i2c_0_csr_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:i2c_0_csr_writedata -> i2c_0:writedata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata       : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest    : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess    : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address        : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read           : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write          : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal mm_interconnect_0_sdram_controller_0_s1_chipselect              : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	signal mm_interconnect_0_sdram_controller_0_s1_readdata                : std_logic_vector(15 downto 0); -- sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	signal mm_interconnect_0_sdram_controller_0_s1_waitrequest             : std_logic;                     -- sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_0_s1_address                 : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	signal mm_interconnect_0_sdram_controller_0_s1_read                    : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_read -> mm_interconnect_0_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_0_s1_byteenable -> mm_interconnect_0_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_0_s1_readdatavalid           : std_logic;                     -- sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_0_s1_write                   : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_write -> mm_interconnect_0_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_sdram_controller_0_s1_writedata               : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	signal mm_interconnect_0_nios_leds_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:nios_leds_s1_chipselect -> nios_leds:chipselect
	signal mm_interconnect_0_nios_leds_s1_readdata                         : std_logic_vector(31 downto 0); -- nios_leds:readdata -> mm_interconnect_0:nios_leds_s1_readdata
	signal mm_interconnect_0_nios_leds_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_leds_s1_address -> nios_leds:address
	signal mm_interconnect_0_nios_leds_s1_write                            : std_logic;                     -- mm_interconnect_0:nios_leds_s1_write -> mm_interconnect_0_nios_leds_s1_write:in
	signal mm_interconnect_0_nios_leds_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_leds_s1_writedata -> nios_leds:writedata
	signal mm_interconnect_0_nios_switches_s1_readdata                     : std_logic_vector(31 downto 0); -- nios_switches:readdata -> mm_interconnect_0:nios_switches_s1_readdata
	signal mm_interconnect_0_nios_switches_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_switches_s1_address -> nios_switches:address
	signal mm_interconnect_0_nios_buttons_s1_readdata                      : std_logic_vector(31 downto 0); -- nios_buttons:readdata -> mm_interconnect_0:nios_buttons_s1_readdata
	signal mm_interconnect_0_nios_buttons_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_buttons_s1_address -> nios_buttons:address
	signal mm_interconnect_0_nios_uartrx_s1_readdata                       : std_logic_vector(31 downto 0); -- nios_uartrx:readdata -> mm_interconnect_0:nios_uartrx_s1_readdata
	signal mm_interconnect_0_nios_uartrx_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_uartrx_s1_address -> nios_uartrx:address
	signal mm_interconnect_0_nios_i2cclk_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:nios_i2cclk_s1_chipselect -> nios_i2cclk:chipselect
	signal mm_interconnect_0_nios_i2cclk_s1_readdata                       : std_logic_vector(31 downto 0); -- nios_i2cclk:readdata -> mm_interconnect_0:nios_i2cclk_s1_readdata
	signal mm_interconnect_0_nios_i2cclk_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_i2cclk_s1_address -> nios_i2cclk:address
	signal mm_interconnect_0_nios_i2cclk_s1_write                          : std_logic;                     -- mm_interconnect_0:nios_i2cclk_s1_write -> mm_interconnect_0_nios_i2cclk_s1_write:in
	signal mm_interconnect_0_nios_i2cclk_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_i2cclk_s1_writedata -> nios_i2cclk:writedata
	signal mm_interconnect_0_nios_uarttx_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:nios_uarttx_s1_chipselect -> nios_uarttx:chipselect
	signal mm_interconnect_0_nios_uarttx_s1_readdata                       : std_logic_vector(31 downto 0); -- nios_uarttx:readdata -> mm_interconnect_0:nios_uarttx_s1_readdata
	signal mm_interconnect_0_nios_uarttx_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_uarttx_s1_address -> nios_uarttx:address
	signal mm_interconnect_0_nios_uarttx_s1_write                          : std_logic;                     -- mm_interconnect_0:nios_uarttx_s1_write -> mm_interconnect_0_nios_uarttx_s1_write:in
	signal mm_interconnect_0_nios_uarttx_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_uarttx_s1_writedata -> nios_uarttx:writedata
	signal mm_interconnect_0_nios_i2cdat_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:nios_i2cdat_s1_chipselect -> nios_i2cdat:chipselect
	signal mm_interconnect_0_nios_i2cdat_s1_readdata                       : std_logic_vector(31 downto 0); -- nios_i2cdat:readdata -> mm_interconnect_0:nios_i2cdat_s1_readdata
	signal mm_interconnect_0_nios_i2cdat_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_i2cdat_s1_address -> nios_i2cdat:address
	signal mm_interconnect_0_nios_i2cdat_s1_write                          : std_logic;                     -- mm_interconnect_0:nios_i2cdat_s1_write -> mm_interconnect_0_nios_i2cdat_s1_write:in
	signal mm_interconnect_0_nios_i2cdat_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_i2cdat_s1_writedata -> nios_i2cdat:writedata
	signal mm_interconnect_0_nios_i2crw_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:nios_i2crw_s1_chipselect -> nios_i2crw:chipselect
	signal mm_interconnect_0_nios_i2crw_s1_readdata                        : std_logic_vector(31 downto 0); -- nios_i2crw:readdata -> mm_interconnect_0:nios_i2crw_s1_readdata
	signal mm_interconnect_0_nios_i2crw_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_i2crw_s1_address -> nios_i2crw:address
	signal mm_interconnect_0_nios_i2crw_s1_write                           : std_logic;                     -- mm_interconnect_0:nios_i2crw_s1_write -> mm_interconnect_0_nios_i2crw_s1_write:in
	signal mm_interconnect_0_nios_i2crw_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_i2crw_s1_writedata -> nios_i2crw:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_nios_7seg_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:nios_7seg_s1_chipselect -> nios_7seg:chipselect
	signal mm_interconnect_0_nios_7seg_s1_readdata                         : std_logic_vector(31 downto 0); -- nios_7seg:readdata -> mm_interconnect_0:nios_7seg_s1_readdata
	signal mm_interconnect_0_nios_7seg_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_7seg_s1_address -> nios_7seg:address
	signal mm_interconnect_0_nios_7seg_s1_write                            : std_logic;                     -- mm_interconnect_0:nios_7seg_s1_write -> mm_interconnect_0_nios_7seg_s1_write:in
	signal mm_interconnect_0_nios_7seg_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_7seg_s1_writedata -> nios_7seg:writedata
	signal mm_interconnect_0_nios_header_conn_s1_chipselect                : std_logic;                     -- mm_interconnect_0:nios_header_conn_s1_chipselect -> nios_header_conn:chipselect
	signal mm_interconnect_0_nios_header_conn_s1_readdata                  : std_logic_vector(31 downto 0); -- nios_header_conn:readdata -> mm_interconnect_0:nios_header_conn_s1_readdata
	signal mm_interconnect_0_nios_header_conn_s1_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_header_conn_s1_address -> nios_header_conn:address
	signal mm_interconnect_0_nios_header_conn_s1_write                     : std_logic;                     -- mm_interconnect_0:nios_header_conn_s1_write -> mm_interconnect_0_nios_header_conn_s1_write:in
	signal mm_interconnect_0_nios_header_conn_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_header_conn_s1_writedata -> nios_header_conn:writedata
	signal mm_interconnect_0_uart_0_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_0_uart_0_s1_readdata                            : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	signal mm_interconnect_0_uart_0_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_0_uart_0_s1_read                                : std_logic;                     -- mm_interconnect_0:uart_0_s1_read -> mm_interconnect_0_uart_0_s1_read:in
	signal mm_interconnect_0_uart_0_s1_begintransfer                       : std_logic;                     -- mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_0_uart_0_s1_write                               : std_logic;                     -- mm_interconnect_0:uart_0_s1_write -> mm_interconnect_0_uart_0_s1_write:in
	signal mm_interconnect_0_uart_0_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	signal mm_interconnect_0_nios_oscdivisor_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:nios_oscdivisor_s1_chipselect -> nios_oscdivisor:chipselect
	signal mm_interconnect_0_nios_oscdivisor_s1_readdata                   : std_logic_vector(31 downto 0); -- nios_oscdivisor:readdata -> mm_interconnect_0:nios_oscdivisor_s1_readdata
	signal mm_interconnect_0_nios_oscdivisor_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_oscdivisor_s1_address -> nios_oscdivisor:address
	signal mm_interconnect_0_nios_oscdivisor_s1_write                      : std_logic;                     -- mm_interconnect_0:nios_oscdivisor_s1_write -> mm_interconnect_0_nios_oscdivisor_s1_write:in
	signal mm_interconnect_0_nios_oscdivisor_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_oscdivisor_s1_writedata -> nios_oscdivisor:writedata
	signal mm_interconnect_0_spi_0_spi_control_port_chipselect             : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	signal mm_interconnect_0_spi_0_spi_control_port_readdata               : std_logic_vector(15 downto 0); -- spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	signal mm_interconnect_0_spi_0_spi_control_port_address                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	signal mm_interconnect_0_spi_0_spi_control_port_read                   : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_read -> mm_interconnect_0_spi_0_spi_control_port_read:in
	signal mm_interconnect_0_spi_0_spi_control_port_write                  : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_write -> mm_interconnect_0_spi_0_spi_control_port_write:in
	signal mm_interconnect_0_spi_0_spi_control_port_writedata              : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	signal nios2_qsys_0_d_irq_irq                                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                   : std_logic_vector(0 downto 0);  -- i2c_0:intr -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                               : std_logic_vector(0 downto 0);  -- jtag_uart_0:av_irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_002_receiver_irq                               : std_logic_vector(0 downto 0);  -- timer_0:irq -> irq_synchronizer_002:receiver_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	signal irq_synchronizer_003_receiver_irq                               : std_logic_vector(0 downto 0);  -- uart_0:irq -> irq_synchronizer_003:receiver_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	signal irq_synchronizer_004_receiver_irq                               : std_logic_vector(0 downto 0);  -- spi_0:irq -> irq_synchronizer_004:receiver_irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal nios2_qsys_0_jtag_debug_module_reset_reset                      : std_logic;                     -- nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                     -- rst_controller_001:reset_req -> [nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [pll_0:rst, pll_1:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_sdram_controller_0_s1_read_ports_inv          : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_read:inv -> sdram_controller_0:az_rd_n
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv    : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_0_s1_byteenable:inv -> sdram_controller_0:az_be_n
	signal mm_interconnect_0_sdram_controller_0_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_write:inv -> sdram_controller_0:az_wr_n
	signal mm_interconnect_0_nios_leds_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_nios_leds_s1_write:inv -> nios_leds:write_n
	signal mm_interconnect_0_nios_i2cclk_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_nios_i2cclk_s1_write:inv -> nios_i2cclk:write_n
	signal mm_interconnect_0_nios_uarttx_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_nios_uarttx_s1_write:inv -> nios_uarttx:write_n
	signal mm_interconnect_0_nios_i2cdat_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_nios_i2cdat_s1_write:inv -> nios_i2cdat:write_n
	signal mm_interconnect_0_nios_i2crw_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_nios_i2crw_s1_write:inv -> nios_i2crw:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_nios_7seg_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_nios_7seg_s1_write:inv -> nios_7seg:write_n
	signal mm_interconnect_0_nios_header_conn_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_nios_header_conn_s1_write:inv -> nios_header_conn:write_n
	signal mm_interconnect_0_uart_0_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_0_uart_0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_uart_0_s1_write:inv -> uart_0:write_n
	signal mm_interconnect_0_nios_oscdivisor_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_nios_oscdivisor_s1_write:inv -> nios_oscdivisor:write_n
	signal mm_interconnect_0_spi_0_spi_control_port_read_ports_inv         : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_read:inv -> spi_0:read_n
	signal mm_interconnect_0_spi_0_spi_control_port_write_ports_inv        : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_write:inv -> spi_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [i2c_0:rst_n, jtag_uart_0:rst_n, nios_7seg:reset_n, nios_buttons:reset_n, nios_header_conn:reset_n, nios_i2cclk:reset_n, nios_i2cdat:reset_n, nios_i2crw:reset_n, nios_leds:reset_n, nios_oscdivisor:reset_n, nios_switches:reset_n, nios_uartrx:reset_n, nios_uarttx:reset_n, spi_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, uart_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [nios2_qsys_0:reset_n, sdram_controller_0:reset_n]

begin

	hps_0 : component nios_hps_system_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			h2f_loan_in               => hps_0_h2f_loan_io_in,               --       h2f_loan_io.in
			h2f_loan_out              => hps_0_h2f_loan_io_out,              --                  .out
			h2f_loan_oe               => hps_0_h2f_loan_io_oe,               --                  .oe
			mem_a                     => hps_0_ddr_mem_a,                    --            memory.mem_a
			mem_ba                    => hps_0_ddr_mem_ba,                   --                  .mem_ba
			mem_ck                    => hps_0_ddr_mem_ck,                   --                  .mem_ck
			mem_ck_n                  => hps_0_ddr_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                   => hps_0_ddr_mem_cke,                  --                  .mem_cke
			mem_cs_n                  => hps_0_ddr_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n                 => hps_0_ddr_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n                 => hps_0_ddr_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                  => hps_0_ddr_mem_we_n,                 --                  .mem_we_n
			mem_reset_n               => hps_0_ddr_mem_reset_n,              --                  .mem_reset_n
			mem_dq                    => hps_0_ddr_mem_dq,                   --                  .mem_dq
			mem_dqs                   => hps_0_ddr_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n                 => hps_0_ddr_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                   => hps_0_ddr_mem_odt,                  --                  .mem_odt
			mem_dm                    => hps_0_ddr_mem_dm,                   --                  .mem_dm
			oct_rzqin                 => hps_0_ddr_oct_rzqin,                --                  .oct_rzqin
			hps_io_sdio_inst_CMD      => hps_0_io_hps_io_sdio_inst_CMD,      --            hps_io.hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0       => hps_0_io_hps_io_sdio_inst_D0,       --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1       => hps_0_io_hps_io_sdio_inst_D1,       --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK      => hps_0_io_hps_io_sdio_inst_CLK,      --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2       => hps_0_io_hps_io_sdio_inst_D2,       --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3       => hps_0_io_hps_io_sdio_inst_D3,       --                  .hps_io_sdio_inst_D3
			hps_io_gpio_inst_LOANIO49 => hps_0_io_hps_io_gpio_inst_LOANIO49, --                  .hps_io_gpio_inst_LOANIO49
			hps_io_gpio_inst_LOANIO50 => hps_0_io_hps_io_gpio_inst_LOANIO50, --                  .hps_io_gpio_inst_LOANIO50
			hps_io_gpio_inst_LOANIO55 => hps_0_io_hps_io_gpio_inst_LOANIO55, --                  .hps_io_gpio_inst_LOANIO55
			hps_io_gpio_inst_LOANIO56 => hps_0_io_hps_io_gpio_inst_LOANIO56, --                  .hps_io_gpio_inst_LOANIO56
			h2f_rst_n                 => open,                               --         h2f_reset.reset_n
			h2f_lw_axi_clk            => pll_0_outclk0_clk,                  --  h2f_lw_axi_clock.clk
			h2f_lw_AWID               => open,                               -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR             => open,                               --                  .awaddr
			h2f_lw_AWLEN              => open,                               --                  .awlen
			h2f_lw_AWSIZE             => open,                               --                  .awsize
			h2f_lw_AWBURST            => open,                               --                  .awburst
			h2f_lw_AWLOCK             => open,                               --                  .awlock
			h2f_lw_AWCACHE            => open,                               --                  .awcache
			h2f_lw_AWPROT             => open,                               --                  .awprot
			h2f_lw_AWVALID            => open,                               --                  .awvalid
			h2f_lw_AWREADY            => open,                               --                  .awready
			h2f_lw_WID                => open,                               --                  .wid
			h2f_lw_WDATA              => open,                               --                  .wdata
			h2f_lw_WSTRB              => open,                               --                  .wstrb
			h2f_lw_WLAST              => open,                               --                  .wlast
			h2f_lw_WVALID             => open,                               --                  .wvalid
			h2f_lw_WREADY             => open,                               --                  .wready
			h2f_lw_BID                => open,                               --                  .bid
			h2f_lw_BRESP              => open,                               --                  .bresp
			h2f_lw_BVALID             => open,                               --                  .bvalid
			h2f_lw_BREADY             => open,                               --                  .bready
			h2f_lw_ARID               => open,                               --                  .arid
			h2f_lw_ARADDR             => open,                               --                  .araddr
			h2f_lw_ARLEN              => open,                               --                  .arlen
			h2f_lw_ARSIZE             => open,                               --                  .arsize
			h2f_lw_ARBURST            => open,                               --                  .arburst
			h2f_lw_ARLOCK             => open,                               --                  .arlock
			h2f_lw_ARCACHE            => open,                               --                  .arcache
			h2f_lw_ARPROT             => open,                               --                  .arprot
			h2f_lw_ARVALID            => open,                               --                  .arvalid
			h2f_lw_ARREADY            => open,                               --                  .arready
			h2f_lw_RID                => open,                               --                  .rid
			h2f_lw_RDATA              => open,                               --                  .rdata
			h2f_lw_RRESP              => open,                               --                  .rresp
			h2f_lw_RLAST              => open,                               --                  .rlast
			h2f_lw_RVALID             => open,                               --                  .rvalid
			h2f_lw_RREADY             => open                                --                  .rready
		);

	i2c_0 : component altera_avalon_i2c
		generic map (
			USE_AV_ST       => 0,
			FIFO_DEPTH      => 4,
			FIFO_DEPTH_LOG2 => 2
		)
		port map (
			clk       => pll_0_outclk0_clk,                        --            clock.clk
			rst_n     => rst_controller_reset_out_reset_ports_inv, --       reset_sink.reset_n
			intr      => irq_synchronizer_receiver_irq(0),         -- interrupt_sender.irq
			addr      => mm_interconnect_0_i2c_0_csr_address,      --              csr.address
			read      => mm_interconnect_0_i2c_0_csr_read,         --                 .read
			write     => mm_interconnect_0_i2c_0_csr_write,        --                 .write
			writedata => mm_interconnect_0_i2c_0_csr_writedata,    --                 .writedata
			readdata  => mm_interconnect_0_i2c_0_csr_readdata,     --                 .readdata
			sda_in    => i2c_peripheral_sda_in,                    --       i2c_serial.sda_in
			scl_in    => i2c_peripheral_scl_in,                    --                 .scl_in
			sda_oe    => i2c_peripheral_sda_oe,                    --                 .sda_oe
			scl_oe    => i2c_peripheral_scl_oe,                    --                 .scl_oe
			src_data  => open,                                     --      (terminated)
			src_valid => open,                                     --      (terminated)
			src_ready => '0',                                      --      (terminated)
			snk_data  => "0000000000000000",                       --      (terminated)
			snk_valid => '0',                                      --      (terminated)
			snk_ready => open                                      --      (terminated)
		);

	jtag_uart_0 : component nios_hps_system_jtag_uart_0
		port map (
			clk            => pll_0_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_001_receiver_irq(0)                             --               irq.irq
		);

	nios2_qsys_0 : component nios_hps_system_nios2_qsys_0
		port map (
			clk                                   => pll_0_outclk1_clk,                                            --                       clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,                 --                   reset_n.reset_n
			reset_req                             => rst_controller_001_reset_out_reset_req,                       --                          .reset_req
			d_address                             => nios2_qsys_0_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                          -- custom_instruction_master.readra
		);

	nios_7seg : component nios_hps_system_nios_7seg
		port map (
			clk        => pll_0_outclk0_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_nios_7seg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_7seg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_7seg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_7seg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_7seg_s1_readdata,        --                    .readdata
			out_port   => nios_7seg_export                                -- external_connection.export
		);

	nios_buttons : component nios_hps_system_nios_buttons
		port map (
			clk      => pll_0_outclk0_clk,                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => mm_interconnect_0_nios_buttons_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_nios_buttons_s1_readdata, --                    .readdata
			in_port  => nios_buttons_export                         -- external_connection.export
		);

	nios_header_conn : component nios_hps_system_nios_header_conn
		port map (
			clk        => pll_0_outclk0_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nios_header_conn_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_header_conn_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_header_conn_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_header_conn_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_header_conn_s1_readdata,        --                    .readdata
			in_port    => nios_header_conn_in_port,                              -- external_connection.export
			out_port   => nios_header_conn_out_port                              --                    .export
		);

	nios_i2cclk : component nios_hps_system_nios_i2cclk
		port map (
			clk        => pll_0_outclk0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_nios_i2cclk_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_i2cclk_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_i2cclk_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_i2cclk_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_i2cclk_s1_readdata,        --                    .readdata
			out_port   => nios_i2cclk_export                                -- external_connection.export
		);

	nios_i2cdat : component nios_hps_system_nios_i2cdat
		port map (
			clk        => pll_0_outclk0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_nios_i2cdat_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_i2cdat_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_i2cdat_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_i2cdat_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_i2cdat_s1_readdata,        --                    .readdata
			in_port    => nios_i2cdat_in_port,                              -- external_connection.export
			out_port   => nios_i2cdat_out_port                              --                    .export
		);

	nios_i2crw : component nios_hps_system_nios_i2cclk
		port map (
			clk        => pll_0_outclk0_clk,                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_nios_i2crw_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_i2crw_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_i2crw_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_i2crw_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_i2crw_s1_readdata,        --                    .readdata
			out_port   => nios_i2crw_export                                -- external_connection.export
		);

	nios_leds : component nios_hps_system_nios_leds
		port map (
			clk        => pll_0_outclk0_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_nios_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_leds_s1_readdata,        --                    .readdata
			out_port   => nios_leds_export                                -- external_connection.export
		);

	nios_oscdivisor : component nios_hps_system_nios_oscdivisor
		port map (
			clk        => pll_0_outclk0_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nios_oscdivisor_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_oscdivisor_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_oscdivisor_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_oscdivisor_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_oscdivisor_s1_readdata,        --                    .readdata
			out_port   => nios_oscdivisor_export                                -- external_connection.export
		);

	nios_switches : component nios_hps_system_nios_switches
		port map (
			clk      => pll_0_outclk0_clk,                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => mm_interconnect_0_nios_switches_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_nios_switches_s1_readdata, --                    .readdata
			in_port  => nios_switches_export                         -- external_connection.export
		);

	nios_uartrx : component nios_hps_system_nios_uartrx
		port map (
			clk      => pll_0_outclk0_clk,                         --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_nios_uartrx_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_nios_uartrx_s1_readdata, --                    .readdata
			in_port  => nios_uartrx_export                         -- external_connection.export
		);

	nios_uarttx : component nios_hps_system_nios_i2cclk
		port map (
			clk        => pll_0_outclk0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_nios_uarttx_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_uarttx_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_uarttx_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_uarttx_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_uarttx_s1_readdata,        --                    .readdata
			out_port   => nios_uarttx_export                                -- external_connection.export
		);

	pll_0 : component nios_hps_system_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			outclk_1 => pll_0_outclk1_clk,       -- outclk1.clk
			outclk_2 => pll_0_sdram_clk,         -- outclk2.clk
			locked   => open                     -- (terminated)
		);

	pll_1 : component nios_hps_system_pll_1
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_1_65_clk,            -- outclk0.clk
			outclk_1 => pll_1_108_clk,           -- outclk1.clk
			outclk_2 => pll_1_86_clk,            -- outclk2.clk
			outclk_3 => pll_1_162_clk,           -- outclk3.clk
			outclk_4 => pll_1_144_clk,           -- outclk4.clk
			locked   => open                     -- (terminated)
		);

	sdram_controller_0 : component nios_hps_system_sdram_controller_0
		port map (
			clk            => pll_0_outclk1_clk,                                            --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                 -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_0_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_0_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_0_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_0_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_0_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_0_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_0_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_0_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_0_wire_we_n                                  --      .export
		);

	spi_0 : component nios_hps_system_spi_0
		port map (
			clk           => pll_0_outclk0_clk,                                        --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                 --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_synchronizer_004_receiver_irq(0),                     --              irq.irq
			MISO          => spi_peripheral_MISO,                                      --         external.export
			MOSI          => spi_peripheral_MOSI,                                      --                 .export
			SCLK          => spi_peripheral_SCLK,                                      --                 .export
			SS_n          => spi_peripheral_SS_n                                       --                 .export
		);

	sysid_qsys_0 : component nios_hps_system_sysid_qsys_0
		port map (
			clock    => pll_0_outclk0_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component nios_hps_system_timer_0
		port map (
			clk        => pll_0_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_002_receiver_irq(0)          --   irq.irq
		);

	uart_0 : component nios_hps_system_uart_0
		port map (
			clk           => pll_0_outclk0_clk,                           --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_0_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_0_s1_readdata,        --                    .readdata
			rxd           => uart_peripheral_rxd,                         -- external_connection.export
			txd           => uart_peripheral_txd,                         --                    .export
			irq           => irq_synchronizer_003_receiver_irq(0)         --                 irq.irq
		);

	mm_interconnect_0 : component nios_hps_system_mm_interconnect_0
		port map (
			pll_0_outclk0_clk                                => pll_0_outclk0_clk,                                            --                              pll_0_outclk0.clk
			pll_0_outclk1_clk                                => pll_0_outclk1_clk,                                            --                              pll_0_outclk1.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset    => rst_controller_reset_out_reset,                               --    jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                           -- nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
			nios2_qsys_0_data_master_address                 => nios2_qsys_0_data_master_address,                             --                   nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest             => nios2_qsys_0_data_master_waitrequest,                         --                                           .waitrequest
			nios2_qsys_0_data_master_byteenable              => nios2_qsys_0_data_master_byteenable,                          --                                           .byteenable
			nios2_qsys_0_data_master_read                    => nios2_qsys_0_data_master_read,                                --                                           .read
			nios2_qsys_0_data_master_readdata                => nios2_qsys_0_data_master_readdata,                            --                                           .readdata
			nios2_qsys_0_data_master_write                   => nios2_qsys_0_data_master_write,                               --                                           .write
			nios2_qsys_0_data_master_writedata               => nios2_qsys_0_data_master_writedata,                           --                                           .writedata
			nios2_qsys_0_data_master_debugaccess             => nios2_qsys_0_data_master_debugaccess,                         --                                           .debugaccess
			nios2_qsys_0_instruction_master_address          => nios2_qsys_0_instruction_master_address,                      --            nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest      => nios2_qsys_0_instruction_master_waitrequest,                  --                                           .waitrequest
			nios2_qsys_0_instruction_master_read             => nios2_qsys_0_instruction_master_read,                         --                                           .read
			nios2_qsys_0_instruction_master_readdata         => nios2_qsys_0_instruction_master_readdata,                     --                                           .readdata
			i2c_0_csr_address                                => mm_interconnect_0_i2c_0_csr_address,                          --                                  i2c_0_csr.address
			i2c_0_csr_write                                  => mm_interconnect_0_i2c_0_csr_write,                            --                                           .write
			i2c_0_csr_read                                   => mm_interconnect_0_i2c_0_csr_read,                             --                                           .read
			i2c_0_csr_readdata                               => mm_interconnect_0_i2c_0_csr_readdata,                         --                                           .readdata
			i2c_0_csr_writedata                              => mm_interconnect_0_i2c_0_csr_writedata,                        --                                           .writedata
			jtag_uart_0_avalon_jtag_slave_address            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,      --              jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,        --                                           .write
			jtag_uart_0_avalon_jtag_slave_read               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,         --                                           .read
			jtag_uart_0_avalon_jtag_slave_readdata           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,     --                                           .readdata
			jtag_uart_0_avalon_jtag_slave_writedata          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,    --                                           .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,  --                                           .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,   --                                           .chipselect
			nios2_qsys_0_jtag_debug_module_address           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --             nios2_qsys_0_jtag_debug_module.address
			nios2_qsys_0_jtag_debug_module_write             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                                           .write
			nios2_qsys_0_jtag_debug_module_read              => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                                           .read
			nios2_qsys_0_jtag_debug_module_readdata          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                                           .readdata
			nios2_qsys_0_jtag_debug_module_writedata         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                                           .writedata
			nios2_qsys_0_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                                           .byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                                           .waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                                           .debugaccess
			nios_7seg_s1_address                             => mm_interconnect_0_nios_7seg_s1_address,                       --                               nios_7seg_s1.address
			nios_7seg_s1_write                               => mm_interconnect_0_nios_7seg_s1_write,                         --                                           .write
			nios_7seg_s1_readdata                            => mm_interconnect_0_nios_7seg_s1_readdata,                      --                                           .readdata
			nios_7seg_s1_writedata                           => mm_interconnect_0_nios_7seg_s1_writedata,                     --                                           .writedata
			nios_7seg_s1_chipselect                          => mm_interconnect_0_nios_7seg_s1_chipselect,                    --                                           .chipselect
			nios_buttons_s1_address                          => mm_interconnect_0_nios_buttons_s1_address,                    --                            nios_buttons_s1.address
			nios_buttons_s1_readdata                         => mm_interconnect_0_nios_buttons_s1_readdata,                   --                                           .readdata
			nios_header_conn_s1_address                      => mm_interconnect_0_nios_header_conn_s1_address,                --                        nios_header_conn_s1.address
			nios_header_conn_s1_write                        => mm_interconnect_0_nios_header_conn_s1_write,                  --                                           .write
			nios_header_conn_s1_readdata                     => mm_interconnect_0_nios_header_conn_s1_readdata,               --                                           .readdata
			nios_header_conn_s1_writedata                    => mm_interconnect_0_nios_header_conn_s1_writedata,              --                                           .writedata
			nios_header_conn_s1_chipselect                   => mm_interconnect_0_nios_header_conn_s1_chipselect,             --                                           .chipselect
			nios_i2cclk_s1_address                           => mm_interconnect_0_nios_i2cclk_s1_address,                     --                             nios_i2cclk_s1.address
			nios_i2cclk_s1_write                             => mm_interconnect_0_nios_i2cclk_s1_write,                       --                                           .write
			nios_i2cclk_s1_readdata                          => mm_interconnect_0_nios_i2cclk_s1_readdata,                    --                                           .readdata
			nios_i2cclk_s1_writedata                         => mm_interconnect_0_nios_i2cclk_s1_writedata,                   --                                           .writedata
			nios_i2cclk_s1_chipselect                        => mm_interconnect_0_nios_i2cclk_s1_chipselect,                  --                                           .chipselect
			nios_i2cdat_s1_address                           => mm_interconnect_0_nios_i2cdat_s1_address,                     --                             nios_i2cdat_s1.address
			nios_i2cdat_s1_write                             => mm_interconnect_0_nios_i2cdat_s1_write,                       --                                           .write
			nios_i2cdat_s1_readdata                          => mm_interconnect_0_nios_i2cdat_s1_readdata,                    --                                           .readdata
			nios_i2cdat_s1_writedata                         => mm_interconnect_0_nios_i2cdat_s1_writedata,                   --                                           .writedata
			nios_i2cdat_s1_chipselect                        => mm_interconnect_0_nios_i2cdat_s1_chipselect,                  --                                           .chipselect
			nios_i2crw_s1_address                            => mm_interconnect_0_nios_i2crw_s1_address,                      --                              nios_i2crw_s1.address
			nios_i2crw_s1_write                              => mm_interconnect_0_nios_i2crw_s1_write,                        --                                           .write
			nios_i2crw_s1_readdata                           => mm_interconnect_0_nios_i2crw_s1_readdata,                     --                                           .readdata
			nios_i2crw_s1_writedata                          => mm_interconnect_0_nios_i2crw_s1_writedata,                    --                                           .writedata
			nios_i2crw_s1_chipselect                         => mm_interconnect_0_nios_i2crw_s1_chipselect,                   --                                           .chipselect
			nios_leds_s1_address                             => mm_interconnect_0_nios_leds_s1_address,                       --                               nios_leds_s1.address
			nios_leds_s1_write                               => mm_interconnect_0_nios_leds_s1_write,                         --                                           .write
			nios_leds_s1_readdata                            => mm_interconnect_0_nios_leds_s1_readdata,                      --                                           .readdata
			nios_leds_s1_writedata                           => mm_interconnect_0_nios_leds_s1_writedata,                     --                                           .writedata
			nios_leds_s1_chipselect                          => mm_interconnect_0_nios_leds_s1_chipselect,                    --                                           .chipselect
			nios_oscdivisor_s1_address                       => mm_interconnect_0_nios_oscdivisor_s1_address,                 --                         nios_oscdivisor_s1.address
			nios_oscdivisor_s1_write                         => mm_interconnect_0_nios_oscdivisor_s1_write,                   --                                           .write
			nios_oscdivisor_s1_readdata                      => mm_interconnect_0_nios_oscdivisor_s1_readdata,                --                                           .readdata
			nios_oscdivisor_s1_writedata                     => mm_interconnect_0_nios_oscdivisor_s1_writedata,               --                                           .writedata
			nios_oscdivisor_s1_chipselect                    => mm_interconnect_0_nios_oscdivisor_s1_chipselect,              --                                           .chipselect
			nios_switches_s1_address                         => mm_interconnect_0_nios_switches_s1_address,                   --                           nios_switches_s1.address
			nios_switches_s1_readdata                        => mm_interconnect_0_nios_switches_s1_readdata,                  --                                           .readdata
			nios_uartrx_s1_address                           => mm_interconnect_0_nios_uartrx_s1_address,                     --                             nios_uartrx_s1.address
			nios_uartrx_s1_readdata                          => mm_interconnect_0_nios_uartrx_s1_readdata,                    --                                           .readdata
			nios_uarttx_s1_address                           => mm_interconnect_0_nios_uarttx_s1_address,                     --                             nios_uarttx_s1.address
			nios_uarttx_s1_write                             => mm_interconnect_0_nios_uarttx_s1_write,                       --                                           .write
			nios_uarttx_s1_readdata                          => mm_interconnect_0_nios_uarttx_s1_readdata,                    --                                           .readdata
			nios_uarttx_s1_writedata                         => mm_interconnect_0_nios_uarttx_s1_writedata,                   --                                           .writedata
			nios_uarttx_s1_chipselect                        => mm_interconnect_0_nios_uarttx_s1_chipselect,                  --                                           .chipselect
			sdram_controller_0_s1_address                    => mm_interconnect_0_sdram_controller_0_s1_address,              --                      sdram_controller_0_s1.address
			sdram_controller_0_s1_write                      => mm_interconnect_0_sdram_controller_0_s1_write,                --                                           .write
			sdram_controller_0_s1_read                       => mm_interconnect_0_sdram_controller_0_s1_read,                 --                                           .read
			sdram_controller_0_s1_readdata                   => mm_interconnect_0_sdram_controller_0_s1_readdata,             --                                           .readdata
			sdram_controller_0_s1_writedata                  => mm_interconnect_0_sdram_controller_0_s1_writedata,            --                                           .writedata
			sdram_controller_0_s1_byteenable                 => mm_interconnect_0_sdram_controller_0_s1_byteenable,           --                                           .byteenable
			sdram_controller_0_s1_readdatavalid              => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --                                           .readdatavalid
			sdram_controller_0_s1_waitrequest                => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --                                           .waitrequest
			sdram_controller_0_s1_chipselect                 => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --                                           .chipselect
			spi_0_spi_control_port_address                   => mm_interconnect_0_spi_0_spi_control_port_address,             --                     spi_0_spi_control_port.address
			spi_0_spi_control_port_write                     => mm_interconnect_0_spi_0_spi_control_port_write,               --                                           .write
			spi_0_spi_control_port_read                      => mm_interconnect_0_spi_0_spi_control_port_read,                --                                           .read
			spi_0_spi_control_port_readdata                  => mm_interconnect_0_spi_0_spi_control_port_readdata,            --                                           .readdata
			spi_0_spi_control_port_writedata                 => mm_interconnect_0_spi_0_spi_control_port_writedata,           --                                           .writedata
			spi_0_spi_control_port_chipselect                => mm_interconnect_0_spi_0_spi_control_port_chipselect,          --                                           .chipselect
			sysid_qsys_0_control_slave_address               => mm_interconnect_0_sysid_qsys_0_control_slave_address,         --                 sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata              => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,        --                                           .readdata
			timer_0_s1_address                               => mm_interconnect_0_timer_0_s1_address,                         --                                 timer_0_s1.address
			timer_0_s1_write                                 => mm_interconnect_0_timer_0_s1_write,                           --                                           .write
			timer_0_s1_readdata                              => mm_interconnect_0_timer_0_s1_readdata,                        --                                           .readdata
			timer_0_s1_writedata                             => mm_interconnect_0_timer_0_s1_writedata,                       --                                           .writedata
			timer_0_s1_chipselect                            => mm_interconnect_0_timer_0_s1_chipselect,                      --                                           .chipselect
			uart_0_s1_address                                => mm_interconnect_0_uart_0_s1_address,                          --                                  uart_0_s1.address
			uart_0_s1_write                                  => mm_interconnect_0_uart_0_s1_write,                            --                                           .write
			uart_0_s1_read                                   => mm_interconnect_0_uart_0_s1_read,                             --                                           .read
			uart_0_s1_readdata                               => mm_interconnect_0_uart_0_s1_readdata,                         --                                           .readdata
			uart_0_s1_writedata                              => mm_interconnect_0_uart_0_s1_writedata,                        --                                           .writedata
			uart_0_s1_begintransfer                          => mm_interconnect_0_uart_0_s1_begintransfer,                    --                                           .begintransfer
			uart_0_s1_chipselect                             => mm_interconnect_0_uart_0_s1_chipselect                        --                                           .chipselect
		);

	irq_mapper : component nios_hps_system_irq_mapper
		port map (
			clk           => pll_0_outclk1_clk,                  --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			sender_irq    => nios2_qsys_0_d_irq_irq              --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	irq_synchronizer_003 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_003_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver3_irq            --             sender.irq
		);

	irq_synchronizer_004 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_004_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver4_irq            --             sender.irq
		);

	rst_controller : component nios_hps_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                          --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_001 : component nios_hps_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => pll_0_outclk1_clk,                          --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_read;

	mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_write;

	mm_interconnect_0_nios_leds_s1_write_ports_inv <= not mm_interconnect_0_nios_leds_s1_write;

	mm_interconnect_0_nios_i2cclk_s1_write_ports_inv <= not mm_interconnect_0_nios_i2cclk_s1_write;

	mm_interconnect_0_nios_uarttx_s1_write_ports_inv <= not mm_interconnect_0_nios_uarttx_s1_write;

	mm_interconnect_0_nios_i2cdat_s1_write_ports_inv <= not mm_interconnect_0_nios_i2cdat_s1_write;

	mm_interconnect_0_nios_i2crw_s1_write_ports_inv <= not mm_interconnect_0_nios_i2crw_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_nios_7seg_s1_write_ports_inv <= not mm_interconnect_0_nios_7seg_s1_write;

	mm_interconnect_0_nios_header_conn_s1_write_ports_inv <= not mm_interconnect_0_nios_header_conn_s1_write;

	mm_interconnect_0_uart_0_s1_read_ports_inv <= not mm_interconnect_0_uart_0_s1_read;

	mm_interconnect_0_uart_0_s1_write_ports_inv <= not mm_interconnect_0_uart_0_s1_write;

	mm_interconnect_0_nios_oscdivisor_s1_write_ports_inv <= not mm_interconnect_0_nios_oscdivisor_s1_write;

	mm_interconnect_0_spi_0_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_read;

	mm_interconnect_0_spi_0_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of nios_hps_system
